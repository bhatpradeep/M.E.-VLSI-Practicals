module inheritence;
parent_class a;
child_class c;
  initial begin
    c = new();
  end
endmodule
