class parent_class;
     bit [31:0] addr;
endclass
 
class child_class extends parent_class;
    bit [31:0] data;
endclass
